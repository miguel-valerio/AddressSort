----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:01:44 04/15/2014 
-- Design Name: 
-- Module Name:    PixelROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- charitional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PixelROM is
	generic(	char_width	:positive := 5;
				line_width	:positive := 4;
				column_width:positive := 3;
				data_width	:positive := 8);
	port(		char			:in std_logic_vector(char_width-1 downto 0);		--selects 1 of the 18 chars
				line			:in std_logic_vector(line_width-1 downto 0);		--selects 1 of the 12 lines
				column		:in std_logic_vector(column_width-1 downto 0);	--selects 1 of the 8 columns
				data			:out std_logic);											--returns 1 pixel
end PixelROM;

architecture Behavioral of PixelROM is

	type ROM is array (0 to 17, 0 to 11) of std_logic_vector (7 downto 0);
	
	constant my_rom: ROM := (
	0 =>(	"00000000",	-- 0
			"01111100",
			"11000110",
			"11001110",
			"11011110",
			"11010110",
			"11110110",
			"11100110",
			"11000110",
			"01111100",
			"00000000",
			"00000000"),
			
	1 =>(	"00000000",	--  1
			"00010000",
			"00110000",
			"11110000",
			"00110000",
			"00110000",
			"00110000",
			"00110000",
			"00110000",
			"11111100",
			"00000000",
			"00000000"),
			
	2 =>(	"00000000",	--  2
			"01111000",
			"11001100",
			"11001100",
			"00001100",
			"00011000",
			"00110000",
			"01100000",
			"11001100",
			"11111100",
			"00000000",
			"00000000"),
			
	3 =>(	"00000000",	--  3
			"01111000",
			"11001100",
			"00001100",
			"00001100",
			"00111000",
			"00001100",
			"00001100",
			"11001100",
			"01111000",
			"00000000",
			"00000000"),
			
	4 =>(	"00000000",	--  4
			"00001100",
			"00011100",
			"00111100",
			"01101100",
			"11001100",
			"11111110",
			"00001100",
			"00001100",
			"00011110",
			"00000000",
			"00000000"),
	
	5 =>(	"00000000",	--  5
			"11111100",
			"11000000",
			"11000000",
			"11000000",
			"11111000",
			"00001100",
			"00001100",
			"11001100",
			"01111000",
			"00000000",
			"00000000"),
			
	6 =>(	"00000000",	--  6
			"00111000",
			"01100000",
			"11000000",
			"11000000",
			"11111000",
			"11001100",
			"11001100",
			"11001100",
			"01111000",
			"00000000",
			"00000000"),
			
	7 =>(	"00000000",	--  7
			"11111110",
			"11000110",
			"11000110",
			"00000110",
			"00001100",
			"00011000",
			"00110000",
			"00110000",
			"00110000",
			"00000000",
			"00000000"),
			
	8 =>(	"00000000",	--  8
			"01111000",
			"11001100",
			"11001100",
			"11101100",
			"01111000",
			"11011100",
			"11001100",
			"11001100",
			"01111000",
			"00000000",
			"00000000"),
			
	9 =>(	"00000000",	--  9
			"01111000",
			"11001100",
			"11001100",
			"11001100",
			"01111100",
			"00011000",
			"00011000",
			"00110000",
			"01110000",
			"00000000",
			"00000000"),
			
	10=>(	"00000000",	--  A
			"00110000",
			"01111000",
			"11001100",
			"11001100",
			"11001100",
			"11111100",
			"11001100",
			"11001100",
			"11001100",
			"00000000",
			"00000000"),
			
	11=>(	"00000000",	--  B
			"11111100",
			"01100110",
			"01100110",
			"01100110",
			"01111100",
			"01100110",
			"01100110",
			"01100110",
			"11111100",
			"00000000",
			"00000000"),
			
	12=>(	"00000000",	--  C
			"00111100",
			"01100110",
			"11000110",
			"11000000",
			"11000000",
			"11000000",
			"11000110",
			"01100110",
			"00111100",
			"00000000",
			"00000000"),
			
	13=>(	"00000000",	--  D
			"11111000",
			"01101100",
			"01100110",
			"01100110",
			"01100110",
			"01100110",
			"01100110",
			"01101100",
			"11111000",
			"00000000",
			"00000000"),
			
	14=>(	"00000000",	--  E
			"11111110",
			"01100010",
			"01100000",
			"01100100",
			"01111100",
			"01100100",
			"01100000",
			"01100010",
			"11111110",
			"00000000",
			"00000000"),
			
	15=>(	"00000000",	--  F
			"11111110",
			"01100110",
			"01100000",
			"01100100",
			"01111100",
			"01100100",
			"01100000",
			"01100000",
			"11110000",
			"00000000",
			"00000000"),
			
	16=>(	"00000000",	--  Space
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000"),
			
	17=>(	"00011000",	--  |
			"00011000",
			"00011000",
			"00011000",
			"00011000",
			"00011000",
			"00011000",
			"00011000",
			"00011000",
			"00011000",
			"00011000",
			"00011000"));

begin

	data <= my_rom (conv_integer(char), conv_integer(line))(conv_integer(column));

end Behavioral;

